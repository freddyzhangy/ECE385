	component lab9_soc is
	end component lab9_soc;

	u0 : component lab9_soc
		port map (
		);

