
module lab9_soc (
	);	

endmodule
