//module timing_controller(	
//									input logic Clk,
//									input logic opener,
//									
//									output logic opener_out
//
//									);
//									
//	always_ff @ (posedge Clk)
//	begin
//	for (int i = 0; i < 200000000; i++);								
//		opener_out = opener;
//	end
//	
//endmodule								